class coverage;




endclass : coverage